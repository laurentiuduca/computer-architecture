`timescale 1ns / 10ps

module capture_20200329_1722_24(clk_of_verifla, la_trigger_matched, SDA, SCL, bitcount, memory_line_id);

output clk_of_verifla;
output la_trigger_matched;
output [32:0] memory_line_id;
output SDA;
output SCL;
output [5:0] bitcount;
reg SDA;
reg SCL;
reg [5:0] bitcount;
reg [32:0] memory_line_id;
reg la_trigger_matched;
reg clk_of_verifla;

parameter PERIOD = 20;
initial    // Clock process for clk_of_verifla
begin
    forever
    begin
        clk_of_verifla = 1'b0;
        #(10); clk_of_verifla = 1'b1;
        #(10);
    end
end

initial begin
#(10);
la_trigger_matched = 0;
memory_line_id=7;
{bitcount,SCL,SDA} = 8'b00000010;
#1310660;
// -------------  Current Time:  1310670*(1ns) 
memory_line_id=0;
{bitcount,SCL,SDA} = 8'b00000010;
#1310660;
// -------------  Current Time:  2621330*(1ns) 
memory_line_id=1;
{bitcount,SCL,SDA} = 8'b00000010;
#1310660;
// -------------  Current Time:  3931990*(1ns) 
memory_line_id=2;
{bitcount,SCL,SDA} = 8'b00000010;
#1310660;
// -------------  Current Time:  5242650*(1ns) 
memory_line_id=3;
{bitcount,SCL,SDA} = 8'b00000010;
#1310660;
// -------------  Current Time:  6553310*(1ns) 
memory_line_id=4;
{bitcount,SCL,SDA} = 8'b00000010;
#1310660;
// -------------  Current Time:  7863970*(1ns) 
memory_line_id=5;
{bitcount,SCL,SDA} = 8'b00000010;
#1310660;
// -------------  Current Time:  9174630*(1ns) 
memory_line_id=6;
{bitcount,SCL,SDA} = 8'b00000010;
#39200;
// -------------  Current Time:  9213830*(1ns) 
memory_line_id=8;
{bitcount,SCL,SDA} = 8'b00000000;
la_trigger_matched = 1;
#9000;
// -------------  Current Time:  9222830*(1ns) 
memory_line_id=9;
{bitcount,SCL,SDA} = 8'b00000001;
#6960;
// -------------  Current Time:  9229790*(1ns) 
memory_line_id=10;
{bitcount,SCL,SDA} = 8'b00000111;
#7940;
// -------------  Current Time:  9237730*(1ns) 
memory_line_id=11;
{bitcount,SCL,SDA} = 8'b00000101;
#7980;
// -------------  Current Time:  9245710*(1ns) 
memory_line_id=12;
{bitcount,SCL,SDA} = 8'b00001011;
#7940;
// -------------  Current Time:  9253650*(1ns) 
memory_line_id=13;
{bitcount,SCL,SDA} = 8'b00001001;
#8000;
// -------------  Current Time:  9261650*(1ns) 
memory_line_id=14;
{bitcount,SCL,SDA} = 8'b00001111;
#7940;
// -------------  Current Time:  9269590*(1ns) 
memory_line_id=15;
{bitcount,SCL,SDA} = 8'b00001101;
#980;
// -------------  Current Time:  9270570*(1ns) 
memory_line_id=16;
{bitcount,SCL,SDA} = 8'b00001100;
#7020;
// -------------  Current Time:  9277590*(1ns) 
memory_line_id=17;
{bitcount,SCL,SDA} = 8'b00010010;
#7920;
// -------------  Current Time:  9285510*(1ns) 
memory_line_id=18;
{bitcount,SCL,SDA} = 8'b00010000;
#8000;
// -------------  Current Time:  9293510*(1ns) 
memory_line_id=19;
{bitcount,SCL,SDA} = 8'b00010110;
#7940;
// -------------  Current Time:  9301450*(1ns) 
memory_line_id=20;
{bitcount,SCL,SDA} = 8'b00010100;
#1020;
// -------------  Current Time:  9302470*(1ns) 
memory_line_id=21;
{bitcount,SCL,SDA} = 8'b00010101;
#6960;
// -------------  Current Time:  9309430*(1ns) 
memory_line_id=22;
{bitcount,SCL,SDA} = 8'b00011011;
#7920;
// -------------  Current Time:  9317350*(1ns) 
memory_line_id=23;
{bitcount,SCL,SDA} = 8'b00011001;
#1000;
// -------------  Current Time:  9318350*(1ns) 
memory_line_id=24;
{bitcount,SCL,SDA} = 8'b00011000;
#7000;
// -------------  Current Time:  9325350*(1ns) 
memory_line_id=25;
{bitcount,SCL,SDA} = 8'b00011110;
#7920;
// -------------  Current Time:  9333270*(1ns) 
memory_line_id=26;
{bitcount,SCL,SDA} = 8'b00011100;
#8000;
// -------------  Current Time:  9341270*(1ns) 
memory_line_id=27;
{bitcount,SCL,SDA} = 8'b00100010;
#7940;
// -------------  Current Time:  9349210*(1ns) 
memory_line_id=28;
{bitcount,SCL,SDA} = 8'b00100000;
#8000;
// -------------  Current Time:  9357210*(1ns) 
memory_line_id=29;
{bitcount,SCL,SDA} = 8'b00100110;
#7920;
// -------------  Current Time:  9365130*(1ns) 
memory_line_id=30;
{bitcount,SCL,SDA} = 8'b00100100;
#320;
// -------------  Current Time:  9365450*(1ns) 
memory_line_id=31;
{bitcount,SCL,SDA} = 8'b00100101;
#680;
// -------------  Current Time:  9366130*(1ns) 
memory_line_id=32;
{bitcount,SCL,SDA} = 8'b00100100;
#7020;
// -------------  Current Time:  9373150*(1ns) 
memory_line_id=33;
{bitcount,SCL,SDA} = 8'b00101010;
#7920;
// -------------  Current Time:  9381070*(1ns) 
memory_line_id=34;
{bitcount,SCL,SDA} = 8'b00101000;
#8000;
// -------------  Current Time:  9389070*(1ns) 
memory_line_id=35;
{bitcount,SCL,SDA} = 8'b00101110;
#7920;
// -------------  Current Time:  9396990*(1ns) 
memory_line_id=36;
{bitcount,SCL,SDA} = 8'b00101100;
#1040;
// -------------  Current Time:  9398030*(1ns) 
memory_line_id=37;
{bitcount,SCL,SDA} = 8'b00101101;
#6960;
// -------------  Current Time:  9404990*(1ns) 
memory_line_id=38;
{bitcount,SCL,SDA} = 8'b00110011;
#7920;
// -------------  Current Time:  9412910*(1ns) 
memory_line_id=39;
{bitcount,SCL,SDA} = 8'b00110001;
#1000;
// -------------  Current Time:  9413910*(1ns) 
memory_line_id=40;
{bitcount,SCL,SDA} = 8'b00110000;
#7000;
// -------------  Current Time:  9420910*(1ns) 
memory_line_id=41;
{bitcount,SCL,SDA} = 8'b00110110;
#7920;
// -------------  Current Time:  9428830*(1ns) 
memory_line_id=42;
{bitcount,SCL,SDA} = 8'b00110100;
#8000;
// -------------  Current Time:  9436830*(1ns) 
memory_line_id=43;
{bitcount,SCL,SDA} = 8'b00111010;
#7920;
// -------------  Current Time:  9444750*(1ns) 
memory_line_id=44;
{bitcount,SCL,SDA} = 8'b00111000;
#1040;
// -------------  Current Time:  9445790*(1ns) 
memory_line_id=45;
{bitcount,SCL,SDA} = 8'b00111001;
#6980;
// -------------  Current Time:  9452770*(1ns) 
memory_line_id=46;
{bitcount,SCL,SDA} = 8'b00111111;
#7920;
// -------------  Current Time:  9460690*(1ns) 
memory_line_id=47;
{bitcount,SCL,SDA} = 8'b00111101;
#1000;
// -------------  Current Time:  9461690*(1ns) 
memory_line_id=48;
{bitcount,SCL,SDA} = 8'b00111100;
#7020;
// -------------  Current Time:  9468710*(1ns) 
memory_line_id=49;
{bitcount,SCL,SDA} = 8'b01000010;
#7920;
// -------------  Current Time:  9476630*(1ns) 
memory_line_id=50;
{bitcount,SCL,SDA} = 8'b01000000;
#1040;
// -------------  Current Time:  9477670*(1ns) 
memory_line_id=51;
{bitcount,SCL,SDA} = 8'b01000001;
#6960;
// -------------  Current Time:  9484630*(1ns) 
memory_line_id=52;
{bitcount,SCL,SDA} = 8'b01000111;
#7920;
// -------------  Current Time:  9492550*(1ns) 
memory_line_id=53;
{bitcount,SCL,SDA} = 8'b01000101;
#280;
// -------------  Current Time:  9492830*(1ns) 
memory_line_id=54;
{bitcount,SCL,SDA} = 8'b01000100;
#7720;
// -------------  Current Time:  9500550*(1ns) 
memory_line_id=55;
{bitcount,SCL,SDA} = 8'b01001010;
#7920;
// -------------  Current Time:  9508470*(1ns) 
memory_line_id=56;
{bitcount,SCL,SDA} = 8'b01001000;
#320;
// -------------  Current Time:  9508790*(1ns) 
memory_line_id=57;
{bitcount,SCL,SDA} = 8'b01001001;
#660;
// -------------  Current Time:  9509450*(1ns) 
memory_line_id=58;
{bitcount,SCL,SDA} = 8'b01001000;
#7020;
// -------------  Current Time:  9516470*(1ns) 
memory_line_id=59;
{bitcount,SCL,SDA} = 8'b01001110;
#7940;
// -------------  Current Time:  9524410*(1ns) 
memory_line_id=60;
{bitcount,SCL,SDA} = 8'b00000011;
#624340;
// -------------  Current Time:  10148750*(1ns) 
memory_line_id=61;
{bitcount,SCL,SDA} = 8'b00000010;
#7960;
// -------------  Current Time:  10156710*(1ns) 
memory_line_id=62;
{bitcount,SCL,SDA} = 8'b00000000;
#9000;
// -------------  Current Time:  10165710*(1ns) 
memory_line_id=63;
{bitcount,SCL,SDA} = 8'b00000001;
#6960;
// -------------  Current Time:  10172670*(1ns) 
memory_line_id=64;
{bitcount,SCL,SDA} = 8'b00000111;
#7920;
// -------------  Current Time:  10180590*(1ns) 
memory_line_id=65;
{bitcount,SCL,SDA} = 8'b00000101;
#8020;
// -------------  Current Time:  10188610*(1ns) 
memory_line_id=66;
{bitcount,SCL,SDA} = 8'b00001011;
#7920;
// -------------  Current Time:  10196530*(1ns) 
memory_line_id=67;
{bitcount,SCL,SDA} = 8'b00001001;
#8000;
// -------------  Current Time:  10204530*(1ns) 
memory_line_id=68;
{bitcount,SCL,SDA} = 8'b00001111;
#7920;
// -------------  Current Time:  10212450*(1ns) 
memory_line_id=69;
{bitcount,SCL,SDA} = 8'b00001101;
#1000;
// -------------  Current Time:  10213450*(1ns) 
memory_line_id=70;
{bitcount,SCL,SDA} = 8'b00001100;
#7000;
// -------------  Current Time:  10220450*(1ns) 
memory_line_id=71;
{bitcount,SCL,SDA} = 8'b00010010;
#7920;
// -------------  Current Time:  10228370*(1ns) 
memory_line_id=72;
{bitcount,SCL,SDA} = 8'b00010000;
#8020;
// -------------  Current Time:  10236390*(1ns) 
memory_line_id=73;
{bitcount,SCL,SDA} = 8'b00010110;
#7900;
// -------------  Current Time:  10244290*(1ns) 
memory_line_id=74;
{bitcount,SCL,SDA} = 8'b00010100;
#1040;
// -------------  Current Time:  10245330*(1ns) 
memory_line_id=75;
{bitcount,SCL,SDA} = 8'b00010101;
#6980;
// -------------  Current Time:  10252310*(1ns) 
memory_line_id=76;
{bitcount,SCL,SDA} = 8'b00011011;
#7920;
// -------------  Current Time:  10260230*(1ns) 
memory_line_id=77;
{bitcount,SCL,SDA} = 8'b00011001;
#980;
// -------------  Current Time:  10261210*(1ns) 
memory_line_id=78;
{bitcount,SCL,SDA} = 8'b00011000;
#7020;
// -------------  Current Time:  10268230*(1ns) 
memory_line_id=79;
{bitcount,SCL,SDA} = 8'b00011110;
#7920;
// -------------  Current Time:  10276150*(1ns) 
memory_line_id=80;
{bitcount,SCL,SDA} = 8'b00011100;
#1040;
// -------------  Current Time:  10277190*(1ns) 
memory_line_id=81;
{bitcount,SCL,SDA} = 8'b00011101;
#6960;
// -------------  Current Time:  10284150*(1ns) 
memory_line_id=82;
{bitcount,SCL,SDA} = 8'b00100011;
#7920;
// -------------  Current Time:  10292070*(1ns) 
memory_line_id=83;
{bitcount,SCL,SDA} = 8'b00100001;
#280;
// -------------  Current Time:  10292350*(1ns) 
memory_line_id=84;
{bitcount,SCL,SDA} = 8'b00100000;
#7740;
// -------------  Current Time:  10300090*(1ns) 
memory_line_id=85;
{bitcount,SCL,SDA} = 8'b00100110;
#7920;
// -------------  Current Time:  10308010*(1ns) 
memory_line_id=86;
{bitcount,SCL,SDA} = 8'b00100100;
#8000;
// -------------  Current Time:  10316010*(1ns) 
memory_line_id=87;
{bitcount,SCL,SDA} = 8'b00101010;
#7920;
// -------------  Current Time:  10323930*(1ns) 
memory_line_id=88;
{bitcount,SCL,SDA} = 8'b00101000;
#8000;
// -------------  Current Time:  10331930*(1ns) 
memory_line_id=89;
{bitcount,SCL,SDA} = 8'b00101110;
#7920;
// -------------  Current Time:  10339850*(1ns) 
memory_line_id=90;
{bitcount,SCL,SDA} = 8'b00101100;
#280;
// -------------  Current Time:  10340130*(1ns) 
memory_line_id=91;
{bitcount,SCL,SDA} = 8'b00101101;
#7720;
// -------------  Current Time:  10347850*(1ns) 
memory_line_id=92;
{bitcount,SCL,SDA} = 8'b00110011;
#7920;
// -------------  Current Time:  10355770*(1ns) 
memory_line_id=93;
{bitcount,SCL,SDA} = 8'b00110001;
#280;
// -------------  Current Time:  10356050*(1ns) 
memory_line_id=94;
{bitcount,SCL,SDA} = 8'b00110000;
#7720;
// -------------  Current Time:  10363770*(1ns) 
memory_line_id=95;
{bitcount,SCL,SDA} = 8'b00110110;
#7920;
// -------------  Current Time:  10371690*(1ns) 
memory_line_id=96;
{bitcount,SCL,SDA} = 8'b00110100;
#8020;
// -------------  Current Time:  10379710*(1ns) 
memory_line_id=97;
{bitcount,SCL,SDA} = 8'b00111010;
#7920;
// -------------  Current Time:  10387630*(1ns) 
memory_line_id=98;
{bitcount,SCL,SDA} = 8'b00111000;
#280;
// -------------  Current Time:  10387910*(1ns) 
memory_line_id=99;
{bitcount,SCL,SDA} = 8'b00111001;
#7720;
// -------------  Current Time:  10395630*(1ns) 
memory_line_id=100;
{bitcount,SCL,SDA} = 8'b00111111;
#7920;
// -------------  Current Time:  10403550*(1ns) 
memory_line_id=101;
{bitcount,SCL,SDA} = 8'b00111101;
#280;
// -------------  Current Time:  10403830*(1ns) 
memory_line_id=102;
{bitcount,SCL,SDA} = 8'b00111100;
#7720;
// -------------  Current Time:  10411550*(1ns) 
memory_line_id=103;
{bitcount,SCL,SDA} = 8'b01000010;
#7920;
// -------------  Current Time:  10419470*(1ns) 
memory_line_id=104;
{bitcount,SCL,SDA} = 8'b01000000;
#280;
// -------------  Current Time:  10419750*(1ns) 
memory_line_id=105;
{bitcount,SCL,SDA} = 8'b01000001;
#7740;
// -------------  Current Time:  10427490*(1ns) 
memory_line_id=106;
{bitcount,SCL,SDA} = 8'b01000111;
#7920;
// -------------  Current Time:  10435410*(1ns) 
memory_line_id=107;
{bitcount,SCL,SDA} = 8'b01000101;
#8000;
// -------------  Current Time:  10443410*(1ns) 
memory_line_id=108;
{bitcount,SCL,SDA} = 8'b01001011;
#7920;
// -------------  Current Time:  10451330*(1ns) 
memory_line_id=109;
{bitcount,SCL,SDA} = 8'b01001001;
#1000;
// -------------  Current Time:  10452330*(1ns) 
memory_line_id=110;
{bitcount,SCL,SDA} = 8'b01001000;
#7000;
// -------------  Current Time:  10459330*(1ns) 
memory_line_id=111;
{bitcount,SCL,SDA} = 8'b01001110;
#7960;
// -------------  Current Time:  10467290*(1ns) 
memory_line_id=112;
{bitcount,SCL,SDA} = 8'b00000011;
#1310660;
// -------------  Current Time:  11777950*(1ns) 
memory_line_id=113;
{bitcount,SCL,SDA} = 8'b00000011;
#1310660;
// -------------  Current Time:  13088610*(1ns) 
memory_line_id=114;
{bitcount,SCL,SDA} = 8'b00000011;
#1310660;
// -------------  Current Time:  14399270*(1ns) 
memory_line_id=115;
{bitcount,SCL,SDA} = 8'b00000011;
#1310660;
// -------------  Current Time:  15709930*(1ns) 
memory_line_id=116;
{bitcount,SCL,SDA} = 8'b00000011;
#1310660;
// -------------  Current Time:  17020590*(1ns) 
memory_line_id=117;
{bitcount,SCL,SDA} = 8'b00000011;
#1310660;
// -------------  Current Time:  18331250*(1ns) 
memory_line_id=118;
{bitcount,SCL,SDA} = 8'b00000011;
#1310660;
// -------------  Current Time:  19641910*(1ns) 
memory_line_id=119;
{bitcount,SCL,SDA} = 8'b00000011;
#1310660;
// -------------  Current Time:  20952570*(1ns) 
memory_line_id=120;
{bitcount,SCL,SDA} = 8'b00000011;
#1310660;
// -------------  Current Time:  22263230*(1ns) 
memory_line_id=121;
{bitcount,SCL,SDA} = 8'b00000011;
#1310660;
// -------------  Current Time:  23573890*(1ns) 
memory_line_id=122;
{bitcount,SCL,SDA} = 8'b00000011;
#1310660;
// -------------  Current Time:  24884550*(1ns) 
memory_line_id=123;
{bitcount,SCL,SDA} = 8'b00000011;
#1310660;
// -------------  Current Time:  26195210*(1ns) 
memory_line_id=124;
{bitcount,SCL,SDA} = 8'b00000011;
#1310660;
// -------------  Current Time:  27505870*(1ns) 
memory_line_id=125;
{bitcount,SCL,SDA} = 8'b00000011;
#1310660;
// -------------  Current Time:  28816530*(1ns) 
memory_line_id=126;
{bitcount,SCL,SDA} = 8'b00000011;
#1310660;
// -------------  Current Time:  30127190*(1ns) 
$finish;
end

initial begin
	$dumpfile("i2c.vcd");
	$dumpvars(0, capture_20200329_1722_24);
end

endmodule
/*
ORIGINAL CAPTURE DUMP
memory_line_id=0: FF FD 02 
memory_line_id=1: FF FD 02 
memory_line_id=2: FF FD 02 
memory_line_id=3: FF FD 02 
memory_line_id=4: FF FD 02 
memory_line_id=5: FF FD 02 
memory_line_id=6: 07 A8 02 
memory_line_id=7: FF FD 02 
memory_line_id=8: 01 C2 00 
memory_line_id=9: 01 5C 01 
memory_line_id=10: 01 8D 07 
memory_line_id=11: 01 8F 05 
memory_line_id=12: 01 8D 0B 
memory_line_id=13: 01 90 09 
memory_line_id=14: 01 8D 0F 
memory_line_id=15: 00 31 0D 
memory_line_id=16: 01 5F 0C 
memory_line_id=17: 01 8C 12 
memory_line_id=18: 01 90 10 
memory_line_id=19: 01 8D 16 
memory_line_id=20: 00 33 14 
memory_line_id=21: 01 5C 15 
memory_line_id=22: 01 8C 1B 
memory_line_id=23: 00 32 19 
memory_line_id=24: 01 5E 18 
memory_line_id=25: 01 8C 1E 
memory_line_id=26: 01 90 1C 
memory_line_id=27: 01 8D 22 
memory_line_id=28: 01 90 20 
memory_line_id=29: 01 8C 26 
memory_line_id=30: 00 10 24 
memory_line_id=31: 00 22 25 
memory_line_id=32: 01 5F 24 
memory_line_id=33: 01 8C 2A 
memory_line_id=34: 01 90 28 
memory_line_id=35: 01 8C 2E 
memory_line_id=36: 00 34 2C 
memory_line_id=37: 01 5C 2D 
memory_line_id=38: 01 8C 33 
memory_line_id=39: 00 32 31 
memory_line_id=40: 01 5E 30 
memory_line_id=41: 01 8C 36 
memory_line_id=42: 01 90 34 
memory_line_id=43: 01 8C 3A 
memory_line_id=44: 00 34 38 
memory_line_id=45: 01 5D 39 
memory_line_id=46: 01 8C 3F 
memory_line_id=47: 00 32 3D 
memory_line_id=48: 01 5F 3C 
memory_line_id=49: 01 8C 42 
memory_line_id=50: 00 34 40 
memory_line_id=51: 01 5C 41 
memory_line_id=52: 01 8C 47 
memory_line_id=53: 00 0E 45 
memory_line_id=54: 01 82 44 
memory_line_id=55: 01 8C 4A 
memory_line_id=56: 00 10 48 
memory_line_id=57: 00 21 49 
memory_line_id=58: 01 5F 48 
memory_line_id=59: 01 8D 4E 
memory_line_id=60: 79 F1 03 
memory_line_id=61: 01 8E 02 
memory_line_id=62: 01 C2 00 
memory_line_id=63: 01 5C 01 
memory_line_id=64: 01 8C 07 
memory_line_id=65: 01 91 05 
memory_line_id=66: 01 8C 0B 
memory_line_id=67: 01 90 09 
memory_line_id=68: 01 8C 0F 
memory_line_id=69: 00 32 0D 
memory_line_id=70: 01 5E 0C 
memory_line_id=71: 01 8C 12 
memory_line_id=72: 01 91 10 
memory_line_id=73: 01 8B 16 
memory_line_id=74: 00 34 14 
memory_line_id=75: 01 5D 15 
memory_line_id=76: 01 8C 1B 
memory_line_id=77: 00 31 19 
memory_line_id=78: 01 5F 18 
memory_line_id=79: 01 8C 1E 
memory_line_id=80: 00 34 1C 
memory_line_id=81: 01 5C 1D 
memory_line_id=82: 01 8C 23 
memory_line_id=83: 00 0E 21 
memory_line_id=84: 01 83 20 
memory_line_id=85: 01 8C 26 
memory_line_id=86: 01 90 24 
memory_line_id=87: 01 8C 2A 
memory_line_id=88: 01 90 28 
memory_line_id=89: 01 8C 2E 
memory_line_id=90: 00 0E 2C 
memory_line_id=91: 01 82 2D 
memory_line_id=92: 01 8C 33 
memory_line_id=93: 00 0E 31 
memory_line_id=94: 01 82 30 
memory_line_id=95: 01 8C 36 
memory_line_id=96: 01 91 34 
memory_line_id=97: 01 8C 3A 
memory_line_id=98: 00 0E 38 
memory_line_id=99: 01 82 39 
memory_line_id=100: 01 8C 3F 
memory_line_id=101: 00 0E 3D 
memory_line_id=102: 01 82 3C 
memory_line_id=103: 01 8C 42 
memory_line_id=104: 00 0E 40 
memory_line_id=105: 01 83 41 
memory_line_id=106: 01 8C 47 
memory_line_id=107: 01 90 45 
memory_line_id=108: 01 8C 4B 
memory_line_id=109: 00 32 49 
memory_line_id=110: 01 5E 48 
memory_line_id=111: 01 8E 4E 
memory_line_id=112: FF FD 03 
memory_line_id=113: FF FD 03 
memory_line_id=114: FF FD 03 
memory_line_id=115: FF FD 03 
memory_line_id=116: FF FD 03 
memory_line_id=117: FF FD 03 
memory_line_id=118: FF FD 03 
memory_line_id=119: FF FD 03 
memory_line_id=120: FF FD 03 
memory_line_id=121: FF FD 03 
memory_line_id=122: FF FD 03 
memory_line_id=123: FF FD 03 
memory_line_id=124: FF FD 03 
memory_line_id=125: FF FD 03 
memory_line_id=126: FF FD 03 
memory_line_id=127: 00 00 06 
*/
